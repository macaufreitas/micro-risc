--------------------------------------------------------------------------------------
---------------- Codigo que implementa o Microprocessador com uma ROM-----------------
--------------------------------------------------------------------------------------

-------- Bibliotecas e Pacotes -------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--------------------------------------

entity MicroprocessadorROM is
	port(
		clk	 : in    std_logic;
		reset  : in    std_logic
	);
end MicroprocessadorROM;

architecture ArquiteturaMicroROM of MicroprocessadorROM is
	--declaração dos sinais
	
	
													
end ArquiteturaMicroROM;